import noc_params::*;

module vc_allocator #(
)(
    input rst,
    input clk,
    input [PORT_NUM-1:0] idle_downstream_vc_i,
    input_block2vc_allocator.vc_allocator ib_if
);

    logic [PORT_NUM-1:0] request_cmd;
    logic [PORT_NUM-1:0] grant;

    logic [PORT_NUM-1:0] is_available_vc, is_available_vc_next;

    separable_input_first_allocator #(
        // .VC_NUM(VC_NUM)
    )
    separable_input_first_allocator (
        .rst(rst),
        .clk(clk),
        .request_i(request_cmd),
        .out_port_i(ib_if.out_port),
        .grant_o(grant)
    );

    /*
    Sequential logic:
    - reset on the rising edge of the rst input;
    - update the availability of downstream Virtual Channels.
    */
    always_ff@(posedge clk, posedge rst)
    begin
        if(rst)
        begin
            is_available_vc <= {PORT_NUM{1'b1}};
        end
        else
        begin
            is_available_vc <= is_available_vc_next;
        end
    end

    /*
    Combinational logic:
    - compute the request matrix for the internal Separable Input-First
      Allocator, by setting to 1 the upstream Virtual Channels which are
      requesting for the allocation of a downstream Virtual Channel and
      whose associated downstream Input Port has at least one available
      Virtual Channel;
    - compute the outputs of the module from the grants matrix obtained
      from the Separable Input-First allocator and update the next
      value for the availability of downstream Virtual Channels if
      they have just been allocated;
    - update the next value for the availability of downstream Virtual
      Channels after their eventual deallocations.
    */
    always_comb
    begin
        is_available_vc_next = is_available_vc;
        for(int up_port = 0; up_port < PORT_NUM; up_port = up_port + 1)
        begin
            // for(int up_vc = 0; up_vc < VC_NUM; up_vc = up_vc + 1)
            // begin
                request_cmd[up_port] = 1'b0;
                ib_if.vc_valid[up_port] = 1'b0;
                // ib_if.vc_new[up_port] = {VC_SIZE{1'bx}};
            // end
        end

        for(int up_port = 0; up_port < PORT_NUM; up_port = up_port + 1)
        begin
            // for(int up_vc = 0; up_vc < VC_NUM; up_vc = up_vc + 1)
            // begin
                if(ib_if.vc_request[up_port] & is_available_vc[ib_if.out_port[up_port]])
                begin
                    request_cmd[up_port] = 1'b1;
                end
            // end
        end

        for(int up_port = 0; up_port < PORT_NUM; up_port = up_port + 1)
        begin
            // for(int up_vc = 0; up_vc < VC_NUM; up_vc = up_vc + 1)
            // begin
                if(grant[up_port])
                begin
                    // ib_if.vc_new[up_port] = assign_downstream_vc(ib_if.out_port[up_port]);
                    ib_if.vc_valid[up_port] = 1'b1;
                    is_available_vc_next[ib_if.out_port[up_port]] = 1'b0;
                end
            // end
        end

        for(int down_port = 0; down_port < PORT_NUM; down_port = down_port + 1)
        begin
            // for(int down_vc = 0; down_vc < VC_NUM; down_vc = down_vc + 1)
            // begin
                if(~is_available_vc[down_port] & idle_downstream_vc_i[down_port])
                begin //! ~is_available_vc[down_port][down_vc] guarantees that 1'b0 set by line 90 is considered.
                    is_available_vc_next[down_port] = 1'b1;
                end
            // end
        end
        
    end

    /*
    Returns the first (starting from 0, without any Round-Robin
    mechanism) Virtual Channel available for allocation from
    the downstream Input Port specified as a parameter.
    */
    //! only 1 VC of only 1 input_port is granted
    // function logic [VC_SIZE-1:0] assign_downstream_vc (input port_t port);
    //     assign_downstream_vc = {VC_SIZE{1'bx}};
    //     // for(int vc = 0; vc < VC_NUM; vc = vc + 1)
    //     // begin
    //         if(is_available_vc[port])
    //         begin
    //             assign_downstream_vc = '0;
    //             break;
    //         end
    //     // end
    // endfunction

endmodule